 /*
 -----------------------------------------------------------------------------
 -- File           : Gray_Nbits_RTL.v
 -----------------------------------------------------------------------------
 */

module gray_Nbits (clk, clk_en, rst, gray_out);
  parameter N = 4;
  parameter SIZE =(N+1);
  parameter Zeros = {SIZE{1'b0}};

  // Place the definition of wires and regs here
  input clk, clk_en, rst;
  output wire [N-1:0] gray_out;
  reg [SIZE-1:0] toogle;
  reg [SIZE-1:0] state;

  reg [N-2:1] or_res;
  integer i;
  integer j;


  // The state of the Gray counter
  always @(posedge clk, negedge rst)
    begin
        if (rst == 1'b0) begin
		    // Initialize state with 1000..00
            state[N] <= 1'b1;
            state[N-1:0] <= 0;
        end
        else begin
		    // Main part of code
            for (j=0; j<(N+1); j=j+1) begin
                if (toogle[j] == 1'b1)
                    state[j] <= ~state[j];
            end
        end
	 end



  // The combinational logic produces the toogle[N:0] signals
  always @(*) begin
        toogle[0] <=  1'b1;
        toogle[1] <= state[0];


        // or_res[i] has the state[i-1:0] bitwise OR
        or_res[1] <= state[0];
        for (i=2; i<N-1; i=i+1) begin
            or_res[i] <= or_res[i-1] | state[i-1];
        end

        for (i=2; i<N; i=i+1) begin
            if ((state[i-1] == 1'b1) && (or_res[i-1] == 1'b0))
                toogle[i] <= 1;
            else
                toogle[i] <= 0;
        end


        if (state[N-2:0] == 0)
            toogle[N] <= 1'b1;
        else
            toogle[N] <= 1'b0;
   end


   assign gray_out = state[N:1];


endmodule
